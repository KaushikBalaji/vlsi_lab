module fibo #parameter(N=32)(
	input clk, rst, 
)
